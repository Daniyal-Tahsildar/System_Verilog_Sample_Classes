class mem_sbd;
    
endclass